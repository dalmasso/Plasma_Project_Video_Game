---------------------------------------------------------------------
-- TITLE: Random Access Memory for Xilinx
-- AUTHOR: Steve Rhoads (rhoadss@yahoo.com)
-- DATE CREATED: 11/06/05
-- FILENAME: ram_xilinx.vhd
-- PROJECT: Plasma CPU core
-- COPYRIGHT: Software placed into the public domain by the author.
--    Software 'as is' without warranty.  Author liable for nothing.
-- DESCRIPTION:
--    Implements the RAM for Spartan 3 Xilinx FPGA
--
--    Compile the MIPS C and assembly code into "test.axf".
--    Run convert.exe to change "test.axf" to "code.txt" which
--    will contain the hex values of the opcodes.
--    Next run "ram_image ram_xilinx.vhd code.txt ram_image.vhd",
--    to create the "ram_image.vhd" file that will have the opcodes
--    correctly placed inside the INIT_00 => strings.
--    Then include ram_image.vhd in the simulation/synthesis.
---------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_misc.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use work.mlite_pack.all;
library UNISIM;
use UNISIM.vcomponents.all;

entity ram is
   generic(memory_type : string := "DEFAULT");
   port(clk               : in std_logic;
        enable            : in std_logic;
        write_byte_enable : in std_logic_vector(3 downto 0);
        address           : in std_logic_vector(31 downto 2);
        data_write        : in std_logic_vector(31 downto 0);
        data_read         : out std_logic_vector(31 downto 0));
end; --entity ram

architecture logic of ram is
begin

   RAMB16_S9_inst0 : RAMB16_S9
   generic map (
INIT_00 => X"afafafafafafafafafafafafafafafaf2308000c241400ac273c243c243c273c",
INIT_01 => X"8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f8f230c008c8c3caf00af00af2340afaf",
INIT_02 => X"acacacac0003373cac038cac8cac8cac8c243c40034040033423038f038f8f8f",
INIT_03 => X"000300ac0300000034038c8c8c8c8c8c8c8c8c8c8c8c3403acacacacacacacac",
INIT_04 => X"248cac1824003c0000038c3c2404242424142c24240424ac00248c243c3c0000",
INIT_05 => X"000003001c24001030008c241430008c24ac0094ac2400183c000003241ca424",
INIT_06 => X"24033c000424a0242410001028300024a0243c0003001030008cac24ac24003c",
INIT_07 => X"102c261026102c001026102c260214002c3a2c3a00000c240200afafafafaf27",
INIT_08 => X"8f028f8f240c240c00142a0000260c0010240c26240c240c001a001600261000",
INIT_09 => X"3c240c3c240c3c240c3c240c3c240c3caf0cafafafafafafafafaf2727038f8f",
INIT_0A => X"0c3c240c3c3c3c3c3c003c3c0c003c240c3c3c1430248c3c1030008c343cac24",
INIT_0B => X"3c240c3c240c3c240c3c240c3c240c3c240c3c240c3c240c3c240c3c240c3c24",
INIT_0C => X"00243c102c26260c000c020c240c3c00000c240c3c020c26102c2600000c240c",
INIT_0D => X"0c270c3c10260c000c000c923c10ae000c020c00000c270c02108e0000008c00",
INIT_0E => X"000c260c3c10021402260c90023c1200000c260c3c100002a210000c020c0000",
INIT_0F => X"0c000c020c02140202269002021200000c260c00103c140226a002000c3c1200",
INIT_10 => X"240c3c3c10260c321402240c000c260c8c02260c0214321200000c260c3c1024",
INIT_11 => X"1400001002260214000c00a002363c24003c3c103c0c003c000c0014343c000c",
INIT_12 => X"03242414002400001000000000000000000000003c1000003c02100200260c00",
INIT_13 => X"008c343c3c1430008c343c2703008f000caf27ac03343cac0000000000343c00",
INIT_14 => X"03008f8f8f00140092260c92240c00140024100092afaf00af270003ac3c1030",
INIT_15 => X"2703008f240caf2727038f8f8f0206260c24341000102c30022400afafaf2727",
INIT_16 => X"3153656c62747267650a0000000000002703008f8c3c10000caf2730038c343c",
INIT_17 => X"796531006e706e724f303030206e6569612020740a00616d20423a0033312030",
INIT_18 => X"37617965613673647475350a62697965340079617965330a7769796532006f61",
INIT_19 => X"0a0a3d6541206820720a3e00616f446f42316f46007539007368380069796561",
INIT_1A => X"00000000000000000000000000000000000037336820660a0d786e6e0a786e75",
INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(31 downto 24),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(31 downto 24),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(3));

   RAMB16_S9_inst1 : RAMB16_S9
   generic map (
INIT_00 => X"b8afaeadacabaaa9a8a7a6a5a4a3a2a1bd000000a560a4a0bd1d8404a5059c1c",
INIT_01 => X"b9b8afaeadacabaaa9a8a7a6a5a4a3a2a1a50086c6c406bb00bb00ba5a1abfb9",
INIT_02 => X"9392919000405a1a06e0a606a606a606a6a50584e0029b401bbd60bb60bbbabf",
INIT_03 => X"00e000c4e0000085a2e09f9d9c9e979695949392919002e09f9d9c9e97969594",
INIT_04 => X"a5a2a2c002a2020582e0420284616303a540c2c6846163404703a24502078000",
INIT_05 => X"0400e000c0c600404200a284404200a2a5a20082a303a2c0020500e084c082c6",
INIT_06 => X"42e00204a1a5c2626200a7406283400540420200e00040420082820282028202",
INIT_07 => X"4042100002404260000240620300606242026303400000134000b0b1b2b3bfbd",
INIT_08 => X"b240b3bf04000400004022501231001200040031040004000020001300100000",
INIT_09 => X"03840004840004840004840004840004b000b1b2b3b4b5b6b7bebfbdbde0b0b1",
INIT_0A => X"00048400041e1715162001060000048400041543420362164042004242026202",
INIT_0B => X"0484000484000484000484000484000484000484000484000484000484000484",
INIT_0C => X"034202406203c400400060008400044000008400040000034042024000008400",
INIT_0D => X"00c4000400c400400000006404007040000000400000c4000000700040006262",
INIT_0E => X"0000a4000400714032310044710440400000a400040000607000400000004000",
INIT_0F => X"0040000000714032023142710040400000a40000000440323162710000044040",
INIT_10 => X"8400040400e4002240320400400031004471e40071402240400000a400040004",
INIT_11 => X"4000004050105040000000509173131200140400060000040000004363030000",
INIT_12 => X"e063634064634000400244024402440244024404040000200191407140310000",
INIT_13 => X"0062630302404200424202bde000bf0000bfbd44e04202624604a48707630300",
INIT_14 => X"e000b0b1bf00400002100004040000510011400002b1bf80b0bd00e044024042",
INIT_15 => X"bde000bf0400bfbdbde0b0b1bf1101100084840000408244111080b0b1bfbdbd",
INIT_16 => X"3265726f6f686f737447000000000000bde000bf4202400000bfbd42e0424202",
INIT_17 => X"206d2e007374752074303078616b206d7262666957007320666f0a003a380031",
INIT_18 => X"2e64206d772e73646f6d2e007974206d2e007464206d2e006f74206d2e007264",
INIT_19 => X"5600207364006569654120007320526d2032702e006d2e0075652e0074206d77",
INIT_1A => X"0000000000000000000000000000000000003834207769430a3e2074433e2065",
INIT_1B => X"0000000000000000000000000000000000000400008024008000000000000000",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(23 downto 16),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(23 downto 16),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(2));

   RAMB16_S9_inst2 : RAMB16_S9
   generic map (
INIT_00 => X"00000000000000000000000000000000ff00000200ff18000f000f000d008d00",
INIT_01 => X"000000000000000000000000000000000000022000002000d800d800ff700000",
INIT_02 => X"0000000000000010000000000000000000010060006060000000000000000000",
INIT_03 => X"0000000000201000000000000000000000000000000000000000000000000000",
INIT_04 => X"00000000002830281000001000ffff0000ff000000ffff001000000d00103020",
INIT_05 => X"20000000ffff00ff000000000000000000000000000028003028000000ff00ff",
INIT_06 => X"0d000021ffff00000000300000003800000d00000000ff000000000000002030",
INIT_07 => X"0000ff00ff00008000ff0000ff200018000000008000020088900000000000ff",
INIT_08 => X"001000000002000200ff009011000291000002ff000200020000000000ff0000",
INIT_09 => X"300b02000b02000b02000b02000b02000000000000000000000000ff00000000",
INIT_0A => X"02000b020000000000f810000028100b02000000ff3c00000000000000200000",
INIT_0B => X"000c02000c02000c02000c02000c02000c02000c02000c02000c02000b02000b",
INIT_0C => X"180d00ff00ff0c02200220000c02009800000c02002002ff0000ff8098020c02",
INIT_0D => X"000c0200ff0c02200200000000ff00200220008000000c022000000000000018",
INIT_0E => X"88000d0200ff10ff100002001000ff9088000d0200ff00f800ff200220008000",
INIT_0F => X"022002200010ff108000001088009080000d0200ff00ff10000018000200ff90",
INIT_10 => X"0d020000ff0d0200ff1000022002000000100d02100000009088000d0200ff00",
INIT_11 => X"000000ff100010000002800010ff007f881000ff00002810200000ff56120000",
INIT_12 => X"00ff00ff1000201800111011101110101011101000ff00f81010ff1080000200",
INIT_13 => X"000000202000000000002000000000000100ff0000002000101020203a002000",
INIT_14 => X"001000000000ff000000020000020000000000000000008000ff10000020ff00",
INIT_15 => X"00000000000200ff000000000010ffff0200000000000000100088000000ff00",
INIT_16 => X"207020616f656d206972000000000000000000000020ff000200ff0000000020",
INIT_17 => X"726f20003a69204d680a303174656c6179696f6e61006866726f0000353a0037",
INIT_18 => X"200a726f20200a72207020007465776f20006520726f20007265776f20006420",
INIT_19 => X"610000736400786e736400006866202066387920007020006d63200065776f20",
INIT_1A => X"0505050508050508070707070606060600003e353169726f002068206f206820",
INIT_1B => X"0000000000000000000000000000000000002000000020080000080505050505",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(15 downto 8),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(15 downto 8),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(1));

   RAMB16_S9_inst3 : RAMB16_S9
   generic map (
INIT_00 => X"4c4844403c3834302c2824201c181410980e006d04fd2a00b800d000b800a801",
INIT_01 => X"504c4844403c3834302c2824201c18141000b82410200060125c1058fc005450",
INIT_02 => X"0c08040000083c0048080c440840043c006000000800000801681360115c5854",
INIT_03 => X"00080c000810121900082c2824201c1814100c08040000082c2824201c181410",
INIT_04 => X"04000007ff2100402108000001feff6304f6080101feff002103009800002525",
INIT_05 => X"40000800effe00fc800000020680000004000000004021140040000802fb00fe",
INIT_06 => X"c0080002f6ff0037300221030a0f250708c000000800fc80000000d000202100",
INIT_07 => X"031ac9149f031a2519bf030ad0252625010d010a2500c50825251014181c20d8",
INIT_08 => X"18251c200a750d7500d2102100017502050875ff207508750008000c00a90f00",
INIT_09 => X"00948600888600848600788600588600108014181c2024282c3034c828081014",
INIT_0A => X"8600ac860000000000090002982500988600000cff1c000010010000500000ff",
INIT_0B => X"00b08600a486009486007c86006886005486003c86002486000c8600f48600dc",
INIT_0C => X"804000be16cff886258625cdec86002500e0d886002575cf130ad02525c5d486",
INIT_0D => X"e0fc8600a0f886258600cd0000a900258625cd2500e0fc86250e000008000021",
INIT_0E => X"25e00c86008121fb2b01750021008a2525e00c86009100090094258625cd2500",
INIT_0F => X"75258625cd21fb2b2101002125082525e00c86007000f92b01002100c5007a25",
INIT_10 => X"20860000401c860ff22b2075258604cd00211c8621040f102525e00c86005a0a",
INIT_11 => X"070000f92a012a0500c0250021ff0fff2500002f02a6250025bf0036783400e0",
INIT_12 => X"08ff01fe2b012525074021402300238023802140001100090021ee2a2501c500",
INIT_13 => X"000020000008020000200018080010002410e800083000002427042580400000",
INIT_14 => X"082510141800f500000175000d750003000a0d000014182510e025080000fc02",
INIT_15 => X"18080010497510e8200810141806f6fc7557300200030a0f061c25101418e020",
INIT_16 => X"32200064742020666e65000000000000180800100000fd00c010e80108002000",
INIT_17 => X"65724d000a6f4f656500303020646967206e726769000a6c6f74000035350000",
INIT_18 => X"520065726d52006561204a00652072724d000a6265724d00642072724d000a77",
INIT_19 => X"6c00002072003e20736400000a6c7444724b2043000a44000a6b43000a72726d",
INIT_1A => X"6c6c6c6cb86c6c0cb4703020f4d0a0940000203632746d6e0000656975006569",
INIT_1B => X"0000000000000000000000000000000000000010102000002070746c6c6c6c6c",
INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DO   => data_read(7 downto 0),
      DOP  => open, 
      ADDR => address(12 downto 2),
      CLK  => clk, 
      DI   => data_write(7 downto 0),
      DIP  => ZERO(0 downto 0),
      EN   => enable,
      SSR  => ZERO(0),
      WE   => write_byte_enable(0));

end; --architecture logic